module MoveGen(
    input logic [8:0] x,
    input logic [8:0] o,
    output logic [8:0] newO);

    logic [8:0] win_play;
    logic [8:0] block_play;
    logic [8:0] fill_play;

                     // row 1
    assign win_play =(o[0] && o[1] && !x[2] && !o[2])? 9'b000_000_100:
                     (o[0] && o[2] && !x[1] && !o[1])? 9'b000_000_010:
                     (o[1] && o[2] && !x[0] && !o[0])? 9'b000_000_001:
                     // row 2
                     (o[3] && o[4] && !x[5] && !o[5])? 9'b000_100_000:
                     (o[3] && o[5] && !x[4] && !o[4])? 9'b000_010_000:
                     (o[4] && o[5] && !x[3] && !o[3])? 9'b000_001_000:
                     // row 3
                     (o[6] && o[7] && !x[8] && !o[8])? 9'b100_000_000:
                     (o[6] && o[8] && !x[7] && !o[7])? 9'b010_000_000:
                     (o[7] && o[8] && !x[6] && !o[6])? 9'b001_000_000:
                     // col 1
                     (o[0] && o[3] && !x[6] && !o[6])? 9'b001_000_000:
                     (o[0] && o[6] && !x[3] && !o[3])? 9'b000_001_000:
                     (o[3] && o[6] && !x[0] && !o[0])? 9'b000_000_001:
                     // col 2
                     (o[1] && o[4] && !x[7] && !o[7])? 9'b010_000_000:
                     (o[1] && o[7] && !x[4] && !o[4])? 9'b000_010_000:
                     (o[4] && o[7] && !x[1] && !o[1])? 9'b000_000_010:
                     // col 3
                     (o[2] && o[5] && !x[8] && !o[8])? 9'b100_000_000:
                     (o[2] && o[8] && !x[5] && !o[5])? 9'b000_100_000:
                     (o[5] && o[8] && !x[2] && !o[2])? 9'b000_000_100:
                     // diag 1
                     (o[0] && o[4] && !x[8] && !o[8])? 9'b100_000_000:
                     (o[0] && o[8] && !x[4] && !o[4])? 9'b000_010_000:
                     (o[4] && o[8] && !x[0] && !o[0])? 9'b000_000_001:
                     // diag 2
                     (o[2] && o[4] && !x[6] && !o[6])? 9'b001_000_000:
                     (o[2] && o[6] && !x[4] && !o[4])? 9'b000_010_000:
                     (o[4] && o[6] && !x[2] && !o[2])? 9'b000_000_100:0;

                        // row 1
    assign block_play = (x[0] && x[1] && !o[2] && !x[2])? 9'b000_000_100:
                        (x[0] && x[2] && !o[1] && !x[1])? 9'b000_000_010:
                        (x[1] && x[2] && !o[0] && !x[0])? 9'b000_000_001:
                        // row 2
                        (x[3] && x[4] && !o[5] && !x[5])? 9'b000_100_000:
                        (x[3] && x[5] && !o[4] && !x[4])? 9'b000_010_000:
                        (x[4] && x[5] && !o[3] && !x[3])? 9'b000_001_000:
                        // row 3
                        (x[6] && x[7] && !o[8] && !x[8])? 9'b100_000_000:
                        (x[6] && x[8] && !o[7] && !x[7])? 9'b010_000_000:
                        (x[7] && x[8] && !o[6] && !x[6])? 9'b001_000_000:
                        // col 1
                        (x[0] && x[3] && !o[6] && !x[6])? 9'b001_000_000:
                        (x[0] && x[6] && !o[3] && !x[3])? 9'b000_001_000:
                        (x[3] && x[6] && !o[0] && !x[0])? 9'b000_000_001:
                        // col 2
                        (x[1] && x[4] && !o[7] && !x[7])? 9'b010_000_000:
                        (x[1] && x[7] && !o[4] && !x[4])? 9'b000_010_000:
                        (x[4] && x[7] && !o[1] && !x[1])? 9'b000_000_010:
                        // col 3
                        (x[2] && x[5] && !o[8] && !x[8])? 9'b100_000_000:
                        (x[2] && x[8] && !o[5] && !x[5])? 9'b000_100_000:
                        (x[5] && x[8] && !o[2] && !x[2])? 9'b000_000_100:
                        // diag 1
                        (x[0] && x[4] && !o[8] && !x[8])? 9'b100_000_000:
                        (x[0] && x[8] && !o[4] && !x[4])? 9'b000_010_000:
                        (x[4] && x[8] && !o[0] && !x[0])? 9'b000_000_001:
                        // diag 2
                        (x[2] && x[4] && !o[6] && !x[6])? 9'b001_000_000:
                        (x[2] && x[6] && !o[4] && !x[4])? 9'b000_010_000:
                        (x[4] && x[6] && !o[2] && !x[2])? 9'b000_000_100:
                        // corners
                        (x[1] && x[3] && !o[0] && !o[2] && !o[6] && !x[0])? 9'b000_000_001:
                        (x[1] && x[5] && !o[0] && !o[2] && !o[8] && !x[2])? 9'b000_000_100:
                        (x[3] && x[7] && !o[0] && !o[6] && !o[8] && !x[6])? 9'b001_000_000:
                        (x[5] && x[7] && !o[2] && !o[6] && !o[8] && !x[8])? 9'b100_000_000:
                        // offset corners
                        (x[1] && x[6] && !o[0] && !o[2] && !o[3] && !x[0])? 9'b000_000_001:
                        (x[2] && x[3] && !o[0] && !o[1] && !o[6] && !x[0])? 9'b000_000_001:
                        (x[0] && x[5] && !o[1] && !o[2] && !o[8] && !x[2])? 9'b000_000_100:
                        (x[1] && x[8] && !o[0] && !o[2] && !o[5] && !x[2])? 9'b000_000_100:
                        (x[0] && x[7] && !o[3] && !o[6] && !o[8] && !x[6])? 9'b001_000_000:
                        (x[3] && x[8] && !o[0] && !o[6] && !o[7] && !x[6])? 9'b001_000_000:
                        (x[5] && x[6] && !o[2] && !o[7] && !o[8] && !x[8])? 9'b100_000_000:
                        (x[2] && x[7] && !o[5] && !o[6] && !o[8] && !x[8])? 9'b100_000_000:0;

    assign fill_play = (!x[0] && !o[0] && x[4])? 9'b000_000_001:
                       (!x[4] && !o[4])? 9'b000_010_000:
                       (!x[1] && !o[1])? 9'b000_000_010:
                       (!x[3] && !o[3])? 9'b000_001_000:
                       (!x[5] && !o[5])? 9'b000_100_000:
                       (!x[7] && !o[7])? 9'b010_000_000:
                       (!x[0] && !o[0])? 9'b000_000_001:                 
                       (!x[2] && !o[2])? 9'b000_000_100:
                       (!x[6] && !o[6])? 9'b001_000_000:
                       (!x[8] && !o[8])? 9'b100_000_000:0;

    logic win;
    logic block;
    logic fill;
    assign win =    | win_play;  
    assign block =  | block_play;
    assign fill =   | fill_play;  

    assign newO = (win)?    o | win_play:
                  (block)?  o | block_play:
                  (fill)?   o | fill_play: o;      
 endmodule